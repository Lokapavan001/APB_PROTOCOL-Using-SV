`ifndef APB_PKG
`define APB_PKG

package apb_pkg;
//`include "interface.sv"
`include "transaction.sv"
`include "generator.sv"
`include "driver.sv"
`include "monitor.sv"
//`include "agent.sv"
`include "predictor.sv"
`include "scoreboard.sv"
`include "environment.sv"
//`include "write_read_test.sv"
//`include "write_test.sv"
//`include "read_test.sv"
`include "random_write_read_test.sv"
`include "slave_error_test.sv"
`include "full_test.sv"
//`include "coverage.sv"

event e1;
endpackage
`endif